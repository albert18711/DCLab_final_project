module Sdram_address (
						RESET_N,
						CLK,
						i_TAKE_FRAME,
						i_640_480_60p,
						i_WR_TO_END,
						i_RE_TO_END,
						o_HEAD_ADDR_1,
						o_MAX_ADDR_1,
						o_HEAD_ADDR_2,
						o_MAX_ADDR_2,
						o_LENGTH
					);

input 

endmodule